# Allocation: Simulator allocated 4685 kB (elbread=427 elab2=4122 kernel=135 sdf=0)
# KERNEL: ASDB file was created in location /home/runner/dataset.asdb
# KERNEL: T=5000 | FLAGS=0000 ANY=0 PULSE=0
# KERNEL: T=15000 | FLAGS=0000 ANY=0 PULSE=0
# KERNEL: T=25000 | FLAGS=0000 ANY=0 PULSE=0
# KERNEL: T=35000 | FLAGS=0000 ANY=0 PULSE=0
# KERNEL: T=45000 | FLAGS=1111 ANY=1 PULSE=1
# KERNEL: T=55000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=65000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=75000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=85000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=95000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=105000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=115000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=125000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=135000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=145000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=155000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=165000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=175000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=185000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=195000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=205000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=215000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=225000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=235000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=245000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=255000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=265000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=275000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=285000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=295000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=305000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=315000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=325000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=335000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=345000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=355000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=365000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=375000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=385000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=395000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=405000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=415000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=425000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=435000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=445000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=455000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=465000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=475000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=485000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=495000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=505000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=515000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=525000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=535000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=545000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=555000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=565000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=575000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=585000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=595000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=605000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=615000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=625000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=635000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=645000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=655000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=665000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=675000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=685000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=695000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=705000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=715000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=725000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=735000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=745000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=755000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=765000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=775000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=785000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=795000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=805000 | FLAGS=1111 ANY=1 PULSE=0
# KERNEL: T=815000 | FLAGS=1111 ANY=1 PULSE=0
# RUNTIME: Info: RUNTIME_0068 testbench.sv (30): $finish called


