// Logic-analyzer style UART RX testbench
`timescale 1ns/1ps

module uart_rx_logic_tb;
    initial begin
        $display("Logic analyzer TB placeholder");
        #1000;
        $finish;
    end
endmodule

